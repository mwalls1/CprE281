module mProj2(F,W,X,Y,Z);
	input W,X,Y,Z;
	output F;
	assign F = (~W&~X&~Y)|(~Y&Z&Z)|(~W&X&Z)|(W&~X&Y&Z);
endmodule
